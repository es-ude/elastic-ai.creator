../../../../vhdl/counter.vhd