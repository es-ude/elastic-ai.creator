library ieee;
use ieee.std_logic_1164.all;


entity $name is
    port (
        $signals
    );
end $name;

architecture rtl of $name is

begin

end rtl;
