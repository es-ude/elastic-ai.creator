../../../../vhdl/padder.vhd