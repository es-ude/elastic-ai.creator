../../../../vhdl/padding_remover.vhd