library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use work.bus_package.all;
    
entity weight_bram is
    generic (
        WEIGHT_NUM : integer := 999;
        BITWIDTH : integer := 8
    );   
    port (
        clk : in std_logic;
        en : in std_logic;
        addr : in std_logic_vector(10-1 downto 0);
        data : out bus_array_4_8
    );
end entity weight_bram;

architecture rtl of weight_bram is
    type weight_bram_array_t is array (0 to WEIGHT_NUM-1) of std_logic_vector(BITWIDTH-1 downto 0);
    signal ROM : weight_bram_array_t := ("00000100","00000000","11111011","11111011","00000011","00001001","00001000","11111101","00000111","11111100","00000110","00000110","11110101","00001001","00001001","00000100","00000010","00000001","00000010","00001001","00000100","00000001","00000000","00000100","00000011","00000000","11111111","00000001","00000011","11111110","11111110","11111000","11111110","11111100","11111110","00000000","11111011","11111100","00000000","11111110","00000011","00000011","11111111","00000000","11111100","00000000","00000011","11111110","11111110","00000011","11111111","00000011","11111100","00000011","11111100","00000100","11111110","00000001","00000000","00000000","00000000","00000000","00000000","11111111","11111110","00000010","11111110","11111111","11110110","11111001","00000000","11110111","11110111","11111111","11111001","11111001","11111010","11111100","00000001","11111011","00000001","00000100","11111101","11111100","00000100","11111100","11111100","11111111","00000101","00000100","11111100","00000000","11111111","11111011","11110110","11110100","11111011","11110110","11111011","00000000","11111011","11111010","00000010","00000010","11111100","00000011","00000000","00000001","00000011","00000000","11111111","00000001","00000100","00000011","00000001","00000011","00001010","00001000","00000101","00001000","00000110","00001011","00000100","00000100","00000011","11111010","00000011","11111011","11111100","11111010","11111011","00000000","11111110","00000101","00000011","00000000","00000010","00000001","11111110","00000011","00000110","11111111","00000100","00000001","11111101","00000101","00000010","00000011","11111011","00000000","11111000","11111001","11111001","11111011","00000000","00000001","00000000","00000110","00000100","00001001","00000111","00000101","00000010","11111111","00000001","11111101","00000010","00000100","00000011","00000000","11111100","00000100","11111100","00000000","00000011","11111011","11111111","00000000","00000001","11111100","00000001","00000011","11111101","11111000","11111111","11111001","11111111","11111100","11111111","11111101","00000011","11111011","00000000","11111111","11111110","00000010","11111101","11111100","00000001","11111100","00000000","11111110","00000101","11111111","00000001","00000001","00000010","00000000","00000000","00000011","00000001","00000100","11111110","00000000","00000101","11111011","11111011","00000011","00000001","11111011","00000011","11111010","00000001","00000000","00000000","00000001","00000101","11111111","11111111","00000000","00000110","00000001","00000011","11111111","00000000","00000101","00000000","00000011","00000010","00000100","00000000","00000100","00000100","11111100","00000011","11111101","11111100","11111000","00000000","11111101","11111111","11111101","00000000","11111011","11111011","11111101","11111001","00000000","00000100","00000110","00001000","00001011","00010101","00010011","00010100","00001011","00010011","00010011","00010011","00001011","00001101","00000110","00000101","00000111","00000101","00000110","00000000","00000001","00000001","11111111","11111100","11111100","00000010","00000101","00000000","11111111","00000101","00000001","11111100","11111101","11111000","11111010","11111001","11111100","11111101","11111001","00000000","11111110","11111101","00000010","00000001","11111110","00000011","11111101","11111100","11111111","00000110","00000001","00000000","00000000","00000010","11111101","11110111","11111110","11110110","11111001","11111101","11111110","00000000","11111111","00000011","00000110","00001010","00000100","00000001","00000001","11111100","00000000","11111011","00000001","00000000","11111110","00000001","11111000","11111000","11111100","11111110","11111100","00000001","00000000","00000001","00000011","00000000","11111110","11111111","11111100","11111010","11111011","11111110","00000010","11111101","11111010","00000010","11111100","00000000","11111111","11111101","00000000","00000011","00000100","11111100","00000001","00000000","00000000","00000101","00000001","00000001","11111110","00000000","00000010","00000000","11111111","11110101","00000000","00000011","11111110","00000001","11111010","00001011","00001101","00000010","00000101","00000001","11111111","00000011","11111111","11111010","11110111","11110001","11110111","11111011","11111101","00000000","00000001","00000001","00001011","00000100","00000110","00001000","00000011","00000001","00000110","00001001","00000001","00000110","00000110","00000110","00000111","00000101","00000011","11111111","11111001","11111110","11111010","00000000","11111110","11111100","00000001","11111100","00000010","11111110","11111110","11111101","00000000","00000011","11111011","11111110","00000010","11111011","11111100","11111011","11111011","11111011","00000100","00000001","11111111","00000010","11111011","00000000","00000001","00000000","00000110","00000000","00000000","00000000","11111111","00000100","00000000","00000101","00000001","00000000","00000001","00000001","11111111","00000000","00000011","00000111","00000110","00000000","00000011","00000101","00000001","00000011","00000010","00000001","00000000","00000011","00000100","00000001","00000000","00001000","00000011","00000110","00000100","00000011","00000110","11111111","00000000","00000011","00000000","00000000","00000110","00000110","00000110","00000110","00000100","00000101","00000110","11111110","00000000","00000100","11111111","11111111","00000011","00000000","11111101","00000011","00000011","11111011","00000011","00000001","11111001","11111100","11111110","00000010","11111010","00000000","00000100","00000101","00000011","00000001","11111110","11111011","11111101","00000000","00000111","00000001","00000000","00000100","11111111","11111111","11111111","00000001","00000001","00000001","11111101","11111110","00000111","00000010","00000111","00000111","11111110","11111100","00000011","00000001","11110111","11111011","00000001","11110111","11111100","11111111","00000110","11111101","11111010","00000010","11111110","11111101","11111010","00000000","11111110","11111010","11111100","11111110","11111101","00000100","00000010","11111101","00000011","11111111","00000101","00000011","00000011","11111110","11111110","00000000","00000111","00000011","11111101","11111100","11111101","00000001","00001000","11111111","00000100","00000001","11111000","00000000","00000011","11111011","11111110","00000100","00000100","00000001","00000101","11111110","00000000","00000000","00000100","00000101","11111110","00000001","00000001","00000011","00000000","00000110","00000001","11111011","00000000","11111011","11111001","11110110","11111111","11111001","11111101","00000001","00000000","11111001","11111001","11111110","11111111","11111110","11111111","11111001","00000000","11111110","00000000","00000010","11111101","00000011","11111011","11111101","00000000","00000001","11111101","11111101","00000000","00000001","11111111","00000000","11111111","11111111","00000001","00000110","00001000","00000000","00000101","00000110","00000100","11111110","11111000","11111101","11111010","00000100","00000100","00000101","11111110","00000011","00000101","00000000","00000000","00000011","00000011","00000111","00000001","00000000","11111110","00000111","00000011","00000000","00000010","00000100","00000011","00001011","00000100","11111101","00000011","11111110","11111101","00000100","00000011","11111011","11111010","11111100","11111101","00000101","00001000","00000010","00000101","11110111","11111100","11111110","00000010","00000001","11110101","11111110","00000001","11111110","00000001","00000000","00000100","11111010","11111111","00000010","11111110","11111101","00000111","00001000","11110111","00000110","00010001","00000001","11111101","00001001","00000001","00001001","00000101","11111001","00000000","00000000","00000011","00001001","00000010","00001110","11111000","00000010","11111011","11111100","00001110","00000011","00000010","11111111","00000100","00000111","11111000","00001000","00000001","11111001","00001010","00000001","00001000","00000110","00000010","11111101","00001010","11111010","11110111","11111101","11110111","00000111","00000101","00000000","11111111","11111010","11111111","11111000","00000111","11111000","00001001","00000111","00000110","11110111","00000010","00000000","11111011","00001000","11111011","00001001","00000101","11110100","00000001","11111111","00000101","11111111","11111101","00000000","11111010","11111110","11111110","00000010","00000100","00000100","00001000","00000000","11111101","11111101","00000110","00000000","00000100","11111010","11111010","11111110","11111101","00001001","11110111","11111110","00001000","11111101","00000010","00000001","11111110","00000011","11111010","00000010","00000101","11111111","00000110","11111011","11110001","00001001","11111011","00000000","00000000","11111110","00000110","00001000","11111001","11111101","00000011","00000001","00000001","00000110","11111111","00000011","00000000","11111111","00001000","00001001","11111010","00000000","11111111","11111011","11111000","00001001","00000101","11111111","11111010","00000001","11110101","11111011","11111111","00000011","11110110","00001000","00000011","00000111","00000000","11111111","00000000","11111011","00001000","00010000","00001001","11111110","00000101","00001001","11111111","11111111","00000111","00000001","11111010","00000100","00000000","00000100","00000001","00000011","00000010","00001000","11111001","11111100","00001011","00000101","11111011","00000011","00000010","00001000","00000101","11111000","00000011","00000000","00000001","00001100","00001000","00001010","00000001","00000011","00000010","00000110","00000001","11111000","00000011","11111011","00000110","00000110","00001010","00000010","11111010","00000011","11110111","11110010","11111011","00001000","11111101","00010001","11111111","11111000","11111010","11111110","11111010","11111110","11110111","11111011","00000101","11111010","00001100","11111111","11110100","11111111","11111100","11111101","11111001","00000000","11111101","11111001","11111010","11111010","00000010","11111011","00000000","00000011","00000001","00001000","11111111","00000001","00000110","00000111","00000101","11111000","00001011","00000011","00001001","11111010","11111111","00000000","00000011","11111001","00000101","00000010","00000110","11111011","11110110","11110110","11111111","00000010","11111001","11111110","00000100","00001000","00000010","11111110","11111100","00000001","00000000","11111000","00000011","00000001","00000001","00000111","11111101","00000000","11110000","11111011","11110100","00000000","00000101","00001010","11110001","11110111","00001010","00000101","11111001","00000111","00010001","11111100","00000000","11111101","00000111","00001011","11110111","00000010","11111000","11111011","00000001","11110110","11111001","00001011","00000000","00001101","11111000","11111011","00001101","11111111","11111110","00001010","00001000","00001110","00001011","11111010","11111001","11111010");
    attribute rom_style : string;
    attribute rom_style of ROM : signal is "auto";
    
    procedure write_and_zero_pad (
        variable addr_w : in integer;
        signal rom : in weight_bram_array_t;
        signal data : out bus_array_4_8
    ) is
    begin
        for ii in 0 to 3 loop
            if addr_w+ii <= WEIGHT_NUM-1 then
                data(ii) <= ROM(addr_w+ii); 
            else
                data(ii) <= (others => '0');
            end if;
        end loop;
    end procedure;
begin
    ROM_process: process(clk)
        variable addr_w : integer;
    begin
        if rising_edge(clk) then
            if (en = '1') then
                addr_w := conv_integer(addr);
                write_and_zero_pad(addr_w, rom, data);
                --data <= bus_array_4_8((ROM(addr_w to addr_w+3)));
            end if;
        end if;
    end process ROM_process;
end architecture rtl;