../../../../vhdl/shift_register.vhd