library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;               -- for type conversions

entity tanh_0 is
    port (
        enable : in std_logic;
        clock  : in std_logic;
        x      : in std_logic_vector(8-1 downto 0);
        y      : out std_logic_vector(8-1 downto 0)
    );
end tanh_0;

architecture rtl of tanh_0 is
    signal signed_x : signed(8-1 downto 0) := (others=>'0');
    signal signed_y : signed(8-1 downto 0) := (others=>'0');
begin
    signed_x <= signed(x);
    y <= std_logic_vector(signed_y);
    tanh_0_process : process(x, signed_x)
    begin
        if signed_x <= -128 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -127 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -126 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -125 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -124 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -123 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -122 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -121 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -120 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -119 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -118 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -117 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -116 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -115 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -114 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -113 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -112 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -111 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -110 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -109 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -108 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -107 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -106 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -105 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -104 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -103 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -102 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -101 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -100 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -99 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -98 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -97 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -96 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -95 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -94 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -93 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -92 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -91 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -90 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -89 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -88 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -87 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -86 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -85 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -84 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -83 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -82 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -81 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -80 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -79 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -78 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -77 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -76 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -75 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -74 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -73 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -72 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -71 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -70 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -69 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -68 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -67 then signed_y <= to_signed(-31, 8);
        elsif signed_x <= -66 then signed_y <= to_signed(-30, 8);
        elsif signed_x <= -65 then signed_y <= to_signed(-30, 8);
        elsif signed_x <= -64 then signed_y <= to_signed(-30, 8);
        elsif signed_x <= -63 then signed_y <= to_signed(-30, 8);
        elsif signed_x <= -62 then signed_y <= to_signed(-30, 8);
        elsif signed_x <= -61 then signed_y <= to_signed(-30, 8);
        elsif signed_x <= -60 then signed_y <= to_signed(-30, 8);
        elsif signed_x <= -59 then signed_y <= to_signed(-30, 8);
        elsif signed_x <= -58 then signed_y <= to_signed(-30, 8);
        elsif signed_x <= -57 then signed_y <= to_signed(-30, 8);
        elsif signed_x <= -56 then signed_y <= to_signed(-30, 8);
        elsif signed_x <= -55 then signed_y <= to_signed(-30, 8);
        elsif signed_x <= -54 then signed_y <= to_signed(-29, 8);
        elsif signed_x <= -53 then signed_y <= to_signed(-29, 8);
        elsif signed_x <= -52 then signed_y <= to_signed(-29, 8);
        elsif signed_x <= -51 then signed_y <= to_signed(-29, 8);
        elsif signed_x <= -50 then signed_y <= to_signed(-29, 8);
        elsif signed_x <= -49 then signed_y <= to_signed(-29, 8);
        elsif signed_x <= -48 then signed_y <= to_signed(-28, 8);
        elsif signed_x <= -47 then signed_y <= to_signed(-28, 8);
        elsif signed_x <= -46 then signed_y <= to_signed(-28, 8);
        elsif signed_x <= -45 then signed_y <= to_signed(-28, 8);
        elsif signed_x <= -44 then signed_y <= to_signed(-28, 8);
        elsif signed_x <= -43 then signed_y <= to_signed(-27, 8);
        elsif signed_x <= -42 then signed_y <= to_signed(-27, 8);
        elsif signed_x <= -41 then signed_y <= to_signed(-27, 8);
        elsif signed_x <= -40 then signed_y <= to_signed(-27, 8);
        elsif signed_x <= -39 then signed_y <= to_signed(-26, 8);
        elsif signed_x <= -38 then signed_y <= to_signed(-26, 8);
        elsif signed_x <= -37 then signed_y <= to_signed(-26, 8);
        elsif signed_x <= -36 then signed_y <= to_signed(-25, 8);
        elsif signed_x <= -35 then signed_y <= to_signed(-25, 8);
        elsif signed_x <= -34 then signed_y <= to_signed(-25, 8);
        elsif signed_x <= -33 then signed_y <= to_signed(-24, 8);
        elsif signed_x <= -32 then signed_y <= to_signed(-24, 8);
        elsif signed_x <= -31 then signed_y <= to_signed(-23, 8);
        elsif signed_x <= -30 then signed_y <= to_signed(-23, 8);
        elsif signed_x <= -29 then signed_y <= to_signed(-23, 8);
        elsif signed_x <= -28 then signed_y <= to_signed(-22, 8);
        elsif signed_x <= -27 then signed_y <= to_signed(-22, 8);
        elsif signed_x <= -26 then signed_y <= to_signed(-21, 8);
        elsif signed_x <= -25 then signed_y <= to_signed(-20, 8);
        elsif signed_x <= -24 then signed_y <= to_signed(-20, 8);
        elsif signed_x <= -23 then signed_y <= to_signed(-19, 8);
        elsif signed_x <= -22 then signed_y <= to_signed(-19, 8);
        elsif signed_x <= -21 then signed_y <= to_signed(-18, 8);
        elsif signed_x <= -20 then signed_y <= to_signed(-17, 8);
        elsif signed_x <= -19 then signed_y <= to_signed(-17, 8);
        elsif signed_x <= -18 then signed_y <= to_signed(-16, 8);
        elsif signed_x <= -17 then signed_y <= to_signed(-15, 8);
        elsif signed_x <= -16 then signed_y <= to_signed(-14, 8);
        elsif signed_x <= -15 then signed_y <= to_signed(-13, 8);
        elsif signed_x <= -14 then signed_y <= to_signed(-13, 8);
        elsif signed_x <= -13 then signed_y <= to_signed(-12, 8);
        elsif signed_x <= -12 then signed_y <= to_signed(-11, 8);
        elsif signed_x <= -11 then signed_y <= to_signed(-10, 8);
        elsif signed_x <= -10 then signed_y <= to_signed(-9, 8);
        elsif signed_x <= -9 then signed_y <= to_signed(-8, 8);
        elsif signed_x <= -8 then signed_y <= to_signed(-7, 8);
        elsif signed_x <= -7 then signed_y <= to_signed(-6, 8);
        elsif signed_x <= -6 then signed_y <= to_signed(-5, 8);
        elsif signed_x <= -5 then signed_y <= to_signed(-4, 8);
        elsif signed_x <= -4 then signed_y <= to_signed(-3, 8);
        elsif signed_x <= -3 then signed_y <= to_signed(-2, 8);
        elsif signed_x <= -2 then signed_y <= to_signed(-1, 8);
        elsif signed_x <= -1 then signed_y <= to_signed(0, 8);
        elsif signed_x <= 0 then signed_y <= to_signed(0, 8);
        elsif signed_x <= 1 then signed_y <= to_signed(0, 8);
        elsif signed_x <= 2 then signed_y <= to_signed(1, 8);
        elsif signed_x <= 3 then signed_y <= to_signed(2, 8);
        elsif signed_x <= 4 then signed_y <= to_signed(3, 8);
        elsif signed_x <= 5 then signed_y <= to_signed(4, 8);
        elsif signed_x <= 6 then signed_y <= to_signed(5, 8);
        elsif signed_x <= 7 then signed_y <= to_signed(6, 8);
        elsif signed_x <= 8 then signed_y <= to_signed(7, 8);
        elsif signed_x <= 9 then signed_y <= to_signed(8, 8);
        elsif signed_x <= 10 then signed_y <= to_signed(9, 8);
        elsif signed_x <= 11 then signed_y <= to_signed(10, 8);
        elsif signed_x <= 12 then signed_y <= to_signed(11, 8);
        elsif signed_x <= 13 then signed_y <= to_signed(12, 8);
        elsif signed_x <= 14 then signed_y <= to_signed(13, 8);
        elsif signed_x <= 15 then signed_y <= to_signed(13, 8);
        elsif signed_x <= 16 then signed_y <= to_signed(14, 8);
        elsif signed_x <= 17 then signed_y <= to_signed(15, 8);
        elsif signed_x <= 18 then signed_y <= to_signed(16, 8);
        elsif signed_x <= 19 then signed_y <= to_signed(17, 8);
        elsif signed_x <= 20 then signed_y <= to_signed(17, 8);
        elsif signed_x <= 21 then signed_y <= to_signed(18, 8);
        elsif signed_x <= 22 then signed_y <= to_signed(19, 8);
        elsif signed_x <= 23 then signed_y <= to_signed(19, 8);
        elsif signed_x <= 24 then signed_y <= to_signed(20, 8);
        elsif signed_x <= 25 then signed_y <= to_signed(20, 8);
        elsif signed_x <= 26 then signed_y <= to_signed(21, 8);
        elsif signed_x <= 27 then signed_y <= to_signed(22, 8);
        elsif signed_x <= 28 then signed_y <= to_signed(22, 8);
        elsif signed_x <= 29 then signed_y <= to_signed(23, 8);
        elsif signed_x <= 30 then signed_y <= to_signed(23, 8);
        elsif signed_x <= 31 then signed_y <= to_signed(23, 8);
        elsif signed_x <= 32 then signed_y <= to_signed(24, 8);
        elsif signed_x <= 33 then signed_y <= to_signed(24, 8);
        elsif signed_x <= 34 then signed_y <= to_signed(25, 8);
        elsif signed_x <= 35 then signed_y <= to_signed(25, 8);
        elsif signed_x <= 36 then signed_y <= to_signed(25, 8);
        elsif signed_x <= 37 then signed_y <= to_signed(26, 8);
        elsif signed_x <= 38 then signed_y <= to_signed(26, 8);
        elsif signed_x <= 39 then signed_y <= to_signed(26, 8);
        elsif signed_x <= 40 then signed_y <= to_signed(27, 8);
        elsif signed_x <= 41 then signed_y <= to_signed(27, 8);
        elsif signed_x <= 42 then signed_y <= to_signed(27, 8);
        elsif signed_x <= 43 then signed_y <= to_signed(27, 8);
        elsif signed_x <= 44 then signed_y <= to_signed(28, 8);
        elsif signed_x <= 45 then signed_y <= to_signed(28, 8);
        elsif signed_x <= 46 then signed_y <= to_signed(28, 8);
        elsif signed_x <= 47 then signed_y <= to_signed(28, 8);
        elsif signed_x <= 48 then signed_y <= to_signed(28, 8);
        elsif signed_x <= 49 then signed_y <= to_signed(29, 8);
        elsif signed_x <= 50 then signed_y <= to_signed(29, 8);
        elsif signed_x <= 51 then signed_y <= to_signed(29, 8);
        elsif signed_x <= 52 then signed_y <= to_signed(29, 8);
        elsif signed_x <= 53 then signed_y <= to_signed(29, 8);
        elsif signed_x <= 54 then signed_y <= to_signed(29, 8);
        elsif signed_x <= 55 then signed_y <= to_signed(30, 8);
        elsif signed_x <= 56 then signed_y <= to_signed(30, 8);
        elsif signed_x <= 57 then signed_y <= to_signed(30, 8);
        elsif signed_x <= 58 then signed_y <= to_signed(30, 8);
        elsif signed_x <= 59 then signed_y <= to_signed(30, 8);
        elsif signed_x <= 60 then signed_y <= to_signed(30, 8);
        elsif signed_x <= 61 then signed_y <= to_signed(30, 8);
        elsif signed_x <= 62 then signed_y <= to_signed(30, 8);
        elsif signed_x <= 63 then signed_y <= to_signed(30, 8);
        elsif signed_x <= 64 then signed_y <= to_signed(30, 8);
        elsif signed_x <= 65 then signed_y <= to_signed(30, 8);
        elsif signed_x <= 66 then signed_y <= to_signed(30, 8);
        elsif signed_x <= 67 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 68 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 69 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 70 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 71 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 72 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 73 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 74 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 75 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 76 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 77 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 78 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 79 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 80 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 81 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 82 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 83 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 84 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 85 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 86 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 87 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 88 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 89 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 90 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 91 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 92 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 93 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 94 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 95 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 96 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 97 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 98 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 99 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 100 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 101 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 102 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 103 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 104 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 105 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 106 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 107 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 108 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 109 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 110 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 111 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 112 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 113 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 114 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 115 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 116 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 117 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 118 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 119 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 120 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 121 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 122 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 123 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 124 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 125 then signed_y <= to_signed(31, 8);
        elsif signed_x <= 126 then signed_y <= to_signed(31, 8);
        else signed_y <= to_signed(31, 8);
        end if;
    end process;
end rtl;
