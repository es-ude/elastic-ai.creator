library ieee;
use ieee.std_logic_1164.all;


entity $name is
    $port
end $name;

architecture rtl of $name is
    $declarations
begin
    $definition
end rtl;
