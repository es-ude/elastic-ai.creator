-- Dummy File for testing implementation of conv1d Design
${total_bits}
${frac_bits}
${in_channels}
${out_channels}
${kernel_size}
${stride}
${padding}
