library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use ieee.std_logic_textio.all;
library ${work_library_name};
use ${work_library_name}.all;
entity ${name}_tb is
    generic (
        DATA_WIDTH : integer := ${data_width};
        THREE_THRESHOLD : integer := ${three_threshold};
        MINUS_THREE_THRESHOLD : integer := ${minus_three_threshold};
        ZERO_OUTPUT : integer := ${zero_output};
        ONE_OUTPUT : integer := ${one_output};
        TMP_THRESHOLD : integer := ${tmp_threshold}
    );
port(
    clk : out std_logic
    );
end entity;
-- architecture rtl of ${name}_tb is
--     constant C_CLK_PERIOD : time := 10 ns;
--     signal clock : std_logic := '0';
--     signal reset : std_logic := '0';
--     signal uut_enable : std_logic := '0';
--     signal x : std_logic_vector(DATA_WIDTH - 1 downto 0);
--     signal y : std_logic_vector(DATA_WIDTH - 1 downto 0);
-- begin
--     CLK_GEN : process
--     begin
--         clock <= '1';
--         wait for C_CLK_PERIOD/2;
--         clock <= '0';
--         wait for C_CLK_PERIOD/2;
--     end process CLK_GEN;
--     RESET_GEN : process
--     begin
--         reset <= '1',
--                 '0' after 20.0*C_CLK_PERIOD;
--     wait;
--     end process RESET_GEN;
--     clk <= clock;
--     test_main : process
--         constant file_inputs:      string := "./data/${name}_q_x.txt";
--         constant file_labels:      string := "./data/${name}_q_y.txt";
--         constant file_pred:      string := "./data/${name}_q_out.txt";
--         file fp_inputs:      text;
--         file fp_labels:      text;
--         file fp_pred:      text;
--         variable line_content:  integer;
--         variable line_num:      line;
--         variable filestatus:    file_open_status;
--         variable input_rd_cnt : integer := 0;
--         variable output_rd_cnt : integer := 0;
--     begin
--         file_open (filestatus, fp_inputs, file_inputs, READ_MODE);
--         report file_inputs & LF & HT & "file_open_status = " &
--                     file_open_status'image(filestatus);
--         assert filestatus = OPEN_OK
--             report "file_open_status /= file_ok"
--             severity FAILURE;
--         file_open (filestatus, fp_labels, file_labels, READ_MODE);
--         report file_labels & LF & HT & "file_open_status = " &
--                     file_open_status'image(filestatus);
--         assert filestatus = OPEN_OK
--             report "file_open_status /= file_ok"
--             severity FAILURE;
--         file_open (filestatus, fp_pred, file_pred, WRITE_MODE);
--         report file_pred & LF & HT & "file_open_status = " &
--                     file_open_status'image(filestatus);
--         assert filestatus = OPEN_OK
--             report "file_open_status /= file_ok"
--             severity FAILURE;
--         uut_enable <= '0';
--         wait until reset='0';
--         wait for C_CLK_PERIOD;
--         uut_enable <= '1';
--         while not ENDFILE (fp_inputs) loop
--             readline (fp_inputs, line_num);
--             read (line_num, line_content);
--             x <= std_logic_vector(to_signed(line_content, DATA_WIDTH));
--             wait for 2*C_CLK_PERIOD;
--             readline (fp_labels, line_num);
--             read (line_num, line_content);
--             report "Correct/Simulated = " & integer'image(line_content) & "/" & integer'image(to_integer(signed(y))) & ", Differece = " & integer'image(line_content - to_integer(signed(y)));
--             write (line_num, to_integer(signed(y)));
--             writeline(fp_pred, line_num);
--         end loop;
--         wait until falling_edge(clock);
--         file_close (fp_inputs);
--         file_close (fp_labels);
--         file_close (fp_pred);
--         report "All files closed.";
--         report "Simulation done.";
--         assert false report "Simulation done. The `assertion failure` is intended to stop this simulation." severity FAILURE;
--     end process ;
--     uut: entity ${work_library_name}.${name}(rtl)
--     port map (
--         enable => uut_enable,
--         clock  => clock,
--         x  => x,
--         y  => y
--     );
-- end architecture;
